** Profile: "SCHEMATIC1-DC"  [ C:\Users\marwa\Desktop\Circ\microphone-SCHEMATIC1-DC.sim ] 

** Creating circuit file "microphone-SCHEMATIC1-DC.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 10 100meg
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\microphone-SCHEMATIC1.net" 


.END
