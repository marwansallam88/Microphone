** Profile: "SCHEMATIC1-time"  [ z:\guc\s6\circuits\project\github\microphone\microphone-schematic1-time.sim ] 

** Creating circuit file "microphone-schematic1-time.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\WINDOWS\pspice.ini file:

*Analysis directives: 
.TRAN  0 100ms 0 1ms 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\microphone-SCHEMATIC1.net" 


.END
